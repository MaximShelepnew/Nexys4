`timescale 1ns / 1ps

`ifndef parameters
`define parameters 

    parameter R = 7;
   // parameter TIMER_BITS = 8;
    parameter FINAL_VALUE = 195;
 
`endif