`timescale 1ns / 1ps

`ifndef parameters
`define parameters 

    parameter D_LENGTH = 5;
 
`endif