//`timescale 1ns / 1ps

//module testbenck_encod;

//wire clk;
//reg ROT_A;
//reg ROT_B;
//reg btn;
//wire [6:0] cathode;

//top_module UUT (clk, ROT_A, ROT_B, btn, cathode);
//assign #10 clk = ~clk;

//integer i = 0;

//initial
//begin
    
//    ROT_A = 0;
//    ROT_B = 0;
//     for (i=0;i<256;i=i+1)
//       // #160 switch = i;
        
//    #10 $finish; 
      
//end

//endmodule
