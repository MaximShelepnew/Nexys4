`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 27.06.2023 21:54:37
// Design Name: 
// Module Name: GREEN
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module GREEN(
    input clk,
    input reset_n,
    input duty,
    input FINAL_VALUE,
    output pwm_out
    );
endmodule
